module tt_um_example (A, B);

    input A;
    output B;

    assign B = A;

endmodule
